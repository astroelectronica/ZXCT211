.title KiCad schematic
.include "C:/AE/ZXCT211/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/ZXCT211/ZXCT211.LIB"
V3 /VSUPPLY 0 DC {VSUPPLY} 
V1 /VIN 0 DC {VIN} 
V2 /VREF 0 DC {VREF} 
R1 /IN- /VIN {RSNS}
XU1 /VREF 0 /VSUPPLY /VIN /IN- /CNV ZXCT211
R2 /CNV /OUT {ROUT}
XU2 /OUT 0 CEU4J2X7R2A103K125AE_s
I1 /IN- 0 DC {ILOAD} 
.end
